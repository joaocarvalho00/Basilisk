`define N_ROWS 4
`define WIDTH 8