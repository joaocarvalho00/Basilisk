`define N_ROWS 			3
`define N_COLUMNS 		3
`define WIDTH 			8
`define ADDR_WIDTH_RAM 	5
`define DEPTH_RAM 		32